`timescale 1ns / 1ps

//////////////////////////////////////////////////////////////////////////////////
// Company: TEC
// Engineer: Carlos Andrey Morales Zamora
// 
// Create Date: 07.03.2025
// Design Name: 
// Module Name: ALU_DUT
// Project Name: LabFPGA2
// 
//////////////////////////////////////////////////////////////////////////////////

module LabFPGA3 #(
	parameter int WIDTH = 24,
	parameter int DIVIDER = 20e6
)(
	input		logic				clk_i,
									rst_i,
									en_reg_i,
									sw_reg_b_i,
									slct_op_i,
	input		logic	[3:0]		cntrl_alu_i,	
	output	logic	[3:0]		flag_o,
	output	logic	[41:0]	display_o,
	output	logic	[1:0]		counter_slct_op_o
						
);
	
	//Internal variables
	logic [WIDTH-1:0] reg_a, reg_b, result, lfsr_a, lfsr_b, signature;
	logic [23:0] display;
	logic [1:0] counter_slct_op;
	logic en_lfsr_a, en_lfsr_b, en_misr;
	
	assign counter_slct_op_o = counter_slct_op;
	
	//Logic select operand
	always_ff @(posedge clk_i) begin
		if(!rst_i) begin counter_slct_op <= 0; end
		else begin
			if(slct_op_i) begin
				if(counter_slct_op == 2) counter_slct_op <= 0;
				else counter_slct_op <= counter_slct_op + 1;
			end
		end
	end
	
	always_comb begin
		case(counter_slct_op) 
			2'b00: display = reg_a;
			2'b01: display = reg_b;
			2'b10: display = signature;
			default: display = 0;
		endcase
	end
	
	//Register logic
	always_ff @(posedge clk_i) begin
		if(!rst_i) begin
			reg_a <= 0;
			reg_b <= 0;
			en_lfsr_a <= 0;
			en_lfsr_b <= 0;
			en_misr <= 0;
		end else begin
			en_lfsr_a <= 0;
			en_lfsr_b <= 0;
			en_misr <= 0;
			if(en_reg_i && counter_slct_op == 2'b00) begin
				reg_a <= lfsr_a;
				en_lfsr_a <= 1;
			end	
			if(en_reg_i && counter_slct_op == 2'b01) begin
				if(!sw_reg_b_i) begin 
					reg_b <= lfsr_b;
					en_lfsr_b <= 1;
				end else reg_b <= result;
			end
			if(en_reg_i && counter_slct_op == 2'b10) begin
				en_misr <= 1;
			end
		end
	end
	
	// Instance for operating A
	LFSR #(
		.WIDTH(WIDTH),
		.POLY(24'hE00201),
		.SEED(24'h2)			// SEED 1
	) LFSR_A (
		.clk_i(clk_i),
		.rst_i(rst_i),
		.en_i(en_lfsr_a),
		.lfsr_o(lfsr_a)
	);

	// Instance for operating B
	LFSR #(
		.WIDTH(WIDTH),
		.POLY(24'hE00201),
		.SEED(24'hABCDE0)		// SEED 2
	) LFSR_B (
		.clk_i(clk_i),
		.rst_i(rst_i),
		.en_i(en_lfsr_b),
		.lfsr_o(lfsr_b)
	);
	
	//MISR to accumulate outputs
	MISR_24bit #(
		 .WIDTH(24),
		 .POLY(24'hE00201)
	) misr (
		 .clk_i(clk_i),
		 .rst_i(rst_i),
		 .en_i(en_misr),
		 .data_i(result),
		 .signature_o(signature)
	);

	ALU_DUT #(
		.WIDTH(WIDTH)
	) ALU (
		.cntrl_alu_i(cntrl_alu_i),
		.reg_a_i(reg_a),
		.reg_b_i(reg_b),
		.flag_o(flag_o),
		.result_o(result)	
	);
	
	seg7_control seg7_crtl (
      .display_i(display),
      .display_o(display_o)
   );
	
endmodule



module ALU_DUT #(
	parameter int WIDTH = 8
)(
	input		logic	[3:0]			cntrl_alu_i,
	input		logic	[WIDTH-1:0]		reg_a_i,
										reg_b_i,
	output		logic	[3:0]			flag_o,
	output		logic	[WIDTH-1:0]		result_o								
);
	
	//Internal variables
	logic	[WIDTH:0] result;
	
	//ALU logic
	always_comb begin
		case(cntrl_alu_i)
			0:	result = reg_a_i + reg_b_i;			//add
			1: result = reg_a_i - reg_b_i;         //sub
			2: result = reg_a_i + 1;            	//increase
			3: result = reg_a_i - 1;					//decrease
			4: result = reg_a_i & reg_b_i;         //and
			5: result = reg_a_i | reg_b_i;        //or
			6: result = ~(reg_a_i);					//not a
			7: result = ~(reg_b_i);						//not b
			8:	result = ~(reg_a_i & reg_b_i);		//nand
			9:	result = reg_a_i ^ reg_b_i;			//xor
			10: result = reg_a_i ~^ reg_b_i;		//xnor
			11: result = reg_a_i << reg_b_i;     	//sll
			12: result = reg_a_i >> reg_b_i;     	//srl   
			13: begin                             	//slt (less than)
					if(reg_a_i < reg_b_i) result = 1;
               else result = 0;
            end
			14: begin                               	//  (greater than or equal to)
               if(reg_b_i <= reg_a_i ) result = 1;
               else result = 0;
               end
         default : result = 'b0;
		endcase
	end
	
	//Flag logic
	always_comb begin
		//flag_o[0] = Z
		flag_o[0] = (result == 0);
		//flag_o[1] = S
		flag_o[1] = result[WIDTH-1];  //1 if negative
		//flag_o[2] = O
		flag_o[2] = result[WIDTH];
		//flag_o[3] = C
		flag_o[3] = result[WIDTH];
	end

	//Output logic
	always_comb begin
		result_o = result[WIDTH-1:0];
	end
	
endmodule

module seg7_control(
    input  logic [23:0] display_i,       
    output logic [41:0] display_o        
);

    logic [6:0] segments [5:0];  // Segments per display

    genvar i;
    generate
        for (i = 0; i < 6; i++) begin : display_gen
            seg7_digit decoder (
                .digit_i    (display_i[i*4 +: 4]),
                .segments_o (segments[i])
            );
        end
    endgenerate

    // Concatenate the 6 groups of 7 bits into a single output vector
    always_comb begin
        display_o = {
            segments[5],
            segments[4],
            segments[3],
            segments[2],
            segments[1],
            segments[0]
        };
    end

endmodule

module seg7_digit(
    input  logic [3:0] digit_i,
    output logic [6:0] segments_o
);

    always_comb begin
        case (digit_i)
			4'h0: segments_o = 7'b100_0000;    //ZERO
			4'h1: segments_o = 7'b111_1001;    //ONE
			4'h2: segments_o = 7'b010_0100;    //TWO
			4'h3: segments_o = 7'b011_0000;    //THREE
			4'h4: segments_o = 7'b001_1001;    //FOUR
			4'h5: segments_o = 7'b001_0010;    //FIVE
			4'h6: segments_o = 7'b000_0010;    //SIX
			4'h7: segments_o = 7'b111_1000;    //SEVEN
			4'h8: segments_o = 7'b000_0000;    //EIGHT
			4'h9: segments_o = 7'b001_1000;    //NINE
			4'ha: segments_o = 7'b000_1000;    //A
			4'hb: segments_o = 7'b000_0011;    //B
			4'hc: segments_o = 7'b100_0110;    //C
			4'hd: segments_o = 7'b010_0001;    //D
			4'he: segments_o = 7'b000_0110;    //E
			4'hf: segments_o = 7'b000_1110;    //F
			default: segments_o = 7'b100_0000;    //ZERO
        endcase
    end

endmodule

module debounce #(
	 parameter int DIVIDER = 20e6
	 )(
    input   logic   clk_i,
                    rst_i,
                    btn_i,
    output  logic   btn_o
 ); 

    logic   [32 : 0]    counter;
    
    logic               start, send;
								
    //Cunter logic
    always_ff @(posedge clk_i) begin
        if(!rst_i) begin
            counter	<= 0;
            start		<= 0;
				send		<= 0;
        end else begin
            if(!btn_i && !start) begin
					start	<= 1;
					send	<= 1;	
				end        
            if(start) begin 
                if(counter  == (DIVIDER - 1)) begin
                    counter <= 0;
                    start   <= 0;           
                end else counter <= counter + 1;
					 send	<= 0;	
            end
        end
	 end
	 
    assign btn_o = send;
    
endmodule


module LFSR #(
    parameter int WIDTH = 8,
    parameter logic [WIDTH-1:0] POLY = 24'hE00201,  // taps (x^24 + x^23 + x^22 + x^17 + 1)
    parameter logic [WIDTH-1:0] SEED = 24'h1
)(
    input	logic 				clk_i,
    input	logic 				rst_i,
	input	logic				en_i,
    output  logic [WIDTH-1:0] 	lfsr_o
);
    logic feedback;

    assign feedback = ^(lfsr_o & POLY);  // XOR of active taps

    always_ff @(posedge clk_i) begin
        if(!rst_i) lfsr_o <= SEED;
        else if(en_i) lfsr_o <= {lfsr_o[WIDTH-2:0], feedback}; 
    end
endmodule

module MISR_24bit #(
    parameter int WIDTH = 24,
    parameter logic [WIDTH-1:0] POLY = 24'hE00201
)(
    input	logic clk_i,
    input  	logic rst_i,
	 input	logic en_i,
    input  	logic [WIDTH-1:0] data_i,
    output 	logic [WIDTH-1:0] signature_o
);

    logic [WIDTH-1:0] misr;
    logic feedback;

    // Calculate XOR feedback of the taps and the MSB bit of the input
    assign feedback = misr[WIDTH-1] ^ data_i[WIDTH-1];

    // XOR Mixture Displacement
    always_ff @(posedge clk_i) begin
        if(!rst_i) misr <= '0;
        else if(en_i) misr <= ({misr[WIDTH-2:0], feedback}) ^ data_i;
    end

    assign signature_o = misr;

endmodule


